module job_q_2.4(
    input  logic [3:0] A,  
    output logic P,D 
);
    assign P = ((!A[3])&(!A[2])&A[1]&(!A[0]))|((!A[3])&(!A[2])&A[1]&A[0])|((!A[3])&A[2]&(!A[1])&A[0])|((!A[3])&A[2]&A[1]&A[0])|(A[3]&(!A[2])&A[1]&A[0])|(A[3]&A[2]&(!A[1])&A[0]);  
    assign D=((!A[3])&(!A[2])&(!A[1])&(!A[0]))|((!A[3])&(!A[2])&A[1]&A[0])|((!A[3])&A[2]&A[1]&(!A[0]))|(A[3]&(!A[2])&(!A[1])&A[0])|(A[3]&A[2]&(!A[1])&(!A[0]))|(A[3]&A[2]&A[1]&A[0]);  

endmodule
